`ifndef ROB
`define ROB
`include "const.v"

module ROB{

}

endmodule
`endif